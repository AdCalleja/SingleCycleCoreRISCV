//! ALU that can perform add, sub, and, or.
//! Additionally output the *result is zero* signal to execute branching control.
module ALU(
    input [31:0]    a,  //! rs1
    input [31:0]    b,  //! rs2 / imm
    input [3:0]     AluCtrl,    //! ALU operation selected from ALU control
    output reg [31:0]   Result,
    output          Zero
    
);

//! Select the operation needed based on AluCtrl, signal generated by ALUControl by decoding instruction.
always@(*) begin : AluOperation
    case(AluCtrl)
        4'b0010: Result = a + b;
        4'b0110: Result = a - b;
        4'b0000: Result = a & b;
        4'b0000: Result = a | b;
        default: Result = 0;
    endcase
end

assign Zero = (Result==0);

endmodule


