//! ALU that can perform add, sub, and, or.
//! Additionally output the *result is zero* signal to execute branching control.
module ALU(
    input [31:0]    a,  //! rs1
    input [31:0]    b,  //! rs2 / imm
    input [3:0]     ALUCtrl,    //! ALU operation selected from ALU control
    output reg [31:0]   Result,
    output          ALUZero
    
);

//! Select the operation needed based on ALUCtrl, signal generated by ALUControl by decoding instruction.
always@(*) begin : AluOperation
    case(ALUCtrl)
        4'b0010: Result = a + b;
        4'b0110: Result = a - b;
        4'b0000: Result = a & b;
        4'b0000: Result = a | b;
        default: Result = 0;
    endcase
end

assign ALUZero = (Result==0);

endmodule


